LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


Entity VideoRamMux is
	Port ( 
	
		-- 68000 signals
		CPUAddress 					: in STD_LOGIC_VECTOR(17 downto 0) ;
		VGAAddress 					: in STD_LOGIC_VECTOR(17 downto 0) ;
		ScrollOffset				: in STD_LOGIC_VECTOR(9 downto 0) ;					-- an offset for scrolling
		VIDEO_RAM_WE_H 			: in STD_LOGIC ;											-- `1`when cpu writes to video ram
		VIDEO_RAM_RE_H 			: in STD_LOGIC ;											-- '1' when cpu reads from video ram
		
		CPU_LDS_L, CPU_UDS_L 	: in std_logic ;											-- low when CPU access one, other or both halves of data bus
				
		-- outputs to the Sram chip
		SRAM_ADDRESS 				: out std_logic_vector(17 downto 0) ;				-- output to address bus of video ram

		SRAM_OE_L 					: out std_logic ;											-- output enable during read and Chip select
		SRAM_CE_L 					: out std_logic ;											-- chip enable to video ram
		SRAM_WE_L 					: out std_logic ;											-- write enable to ram when CPU writes otherwise read
		SRAM_LB_L 					: out std_logic ;											-- byte enable signals for lower half of data bus note CPU only writes to one half not the other
		SRAM_UB_L 					: out std_logic ; 										-- byte enable signals for lower half of data bus note CPU only writes to one half not the other
		
		-- graphics chip signals
		GraphicsAddress			: in Std_logic_Vector(17 downto 0) ;
		GraphicsUDS_L				: in Std_logic ;
		GraphicsLDS_L				: in Std_logic ;
		GraphicsRW					: in Std_logic ;
		GraphicsCE_L				: in Std_logic ;
		GraphicsOE_L				: in Std_logic;
		GraphicsBusy_H				: in Std_logic
);	
end;

Architecture a of VideoRamMux is
begin
	process(CPUAddress, VGAAddress, VIDEO_RAM_WE_H, VIDEO_RAM_RE_H, CPU_LDS_L, CPU_UDS_L, GraphicsBusy_H, GraphicsAddress, GraphicsOE_L, GraphicsCE_L, GraphicsRW, GraphicsUDS_L, GraphicsLDS_L, ScrollOffset)
	begin
	
		-- default signals assume the VGA display controller is always accessing Ram
		
		SRAM_ADDRESS 	<= VGAAddress ;
		SRAM_OE_L 		<= '0' ;
		SRAM_CE_L 		<= '0' ;
		SRAM_WE_L 		<= '1' ;															-- read only
		SRAM_LB_L 		<= '0' ;															-- select both halves of the data bus even though only 1 half is used
		SRAM_UB_L 		<= '0' ;

		-- if the graphics controller wants access to the sram
		-- then switch over the mux to present graphics controller signal to the Sram
		
		If(GraphicsBusy_H = '1')	then												-- graphics controller accessing Ram
			SRAM_ADDRESS(17 downto 9) 	<= ScrollOffset(8 downto 0) + GraphicsAddress(17 downto 9) ;		-- add the offset for scrolling
			SRAM_ADDRESS(8 downto 0) 	<= GraphicsAddress(8 downto 0) ;
			SRAM_OE_L 						<= GraphicsOE_L ;
			SRAM_CE_L 						<= GraphicsCE_L ;
			SRAM_WE_L 						<= GraphicsRW ;								-- read only
			SRAM_LB_L 						<= GraphicsLDS_L ;							-- select both halves of the data bus even though only 1 half is used
			SRAM_UB_L 						<= GraphicsUDS_L ;
			
		elsif((VIDEO_RAM_RE_H = '1' or VIDEO_RAM_WE_H = '1')) then		-- if CPU accessing video ram
			SRAM_ADDRESS(17 downto 9) 	<= ScrollOffset(8 downto 0) + CPUAddress(17 downto 9) ;		-- add the offset for scrolling
			SRAM_ADDRESS(8 downto 0) 	<= CPUAddress(8 downto 0) ;
			
			-- switch the video ram over to take signals driven from CPU in place of VGA controller
			SRAM_LB_L 			<= CPU_LDS_L ;
			SRAM_UB_L 			<= CPU_UDS_L ;
			
			if(VIDEO_RAM_RE_H = '1') then										-- if CPU reading from video ram
				SRAM_CE_L 		<= '0';			
				SRAM_OE_L 		<= '0' ;		
				SRAM_WE_L 		<= '1' ;
			elsif(VIDEO_RAM_WE_H = '1')	then								-- if CPU writing to video ram
				SRAM_CE_L 		<= '0';
				SRAM_OE_L 		<= '1' ;
 			SRAM_WE_L 		<= '0' ;	
			end if;
		end if ;
	end process ;
end a ;
